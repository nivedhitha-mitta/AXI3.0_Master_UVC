parameter ADDR_WIDTH = 8;//32;
parameter DATA_WIDTH = 128;